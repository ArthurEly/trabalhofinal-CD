library verilog;
use verilog.vl_types.all;
entity controlevisor_vlg_vec_tst is
end controlevisor_vlg_vec_tst;
