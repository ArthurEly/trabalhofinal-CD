library verilog;
use verilog.vl_types.all;
entity REG_1BIT_vlg_vec_tst is
end REG_1BIT_vlg_vec_tst;
