library verilog;
use verilog.vl_types.all;
entity mux16busx1_vlg_vec_tst is
end mux16busx1_vlg_vec_tst;
