library verilog;
use verilog.vl_types.all;
entity display_utils is
    port(
        a               : out    vl_logic;
        in_e            : in     vl_logic;
        d0              : in     vl_logic;
        b               : out    vl_logic;
        in_2            : in     vl_logic;
        in_d            : in     vl_logic;
        c               : out    vl_logic;
        in_n            : in     vl_logic;
        in_o            : in     vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        in_1            : in     vl_logic;
        g               : out    vl_logic
    );
end display_utils;
