library verilog;
use verilog.vl_types.all;
entity display_utils_vlg_vec_tst is
end display_utils_vlg_vec_tst;
