library verilog;
use verilog.vl_types.all;
entity \trabalhofinalfinal__vlg_sample_tst\ is
    port(
        clock           : in     vl_logic;
        confirma_DA     : in     vl_logic;
        confirma_funcao : in     vl_logic;
        sw0             : in     vl_logic;
        sw1             : in     vl_logic;
        sw2             : in     vl_logic;
        sw3             : in     vl_logic;
        sw4             : in     vl_logic;
        sw5             : in     vl_logic;
        sw6             : in     vl_logic;
        sw7             : in     vl_logic;
        sw8             : in     vl_logic;
        sw9             : in     vl_logic;
        troca_funcao    : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end \trabalhofinalfinal__vlg_sample_tst\;
