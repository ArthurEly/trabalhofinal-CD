library verilog;
use verilog.vl_types.all;
entity MAQUINA_A_vlg_vec_tst is
end MAQUINA_A_vlg_vec_tst;
