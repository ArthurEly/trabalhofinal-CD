library verilog;
use verilog.vl_types.all;
entity MAQUINA_C_vlg_vec_tst is
end MAQUINA_C_vlg_vec_tst;
