library verilog;
use verilog.vl_types.all;
entity MEM_16ADD_SWAP_vlg_vec_tst is
end MEM_16ADD_SWAP_vlg_vec_tst;
