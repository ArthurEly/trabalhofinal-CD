library verilog;
use verilog.vl_types.all;
entity REG_1BYTE_SWAP_vlg_vec_tst is
end REG_1BYTE_SWAP_vlg_vec_tst;
