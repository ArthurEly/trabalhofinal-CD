library verilog;
use verilog.vl_types.all;
entity MAQUINA_B_vlg_vec_tst is
end MAQUINA_B_vlg_vec_tst;
