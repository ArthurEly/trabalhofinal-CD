library verilog;
use verilog.vl_types.all;
entity trabalhofinal_swap_vlg_vec_tst is
end trabalhofinal_swap_vlg_vec_tst;
