library verilog;
use verilog.vl_types.all;
entity decoddisplay_vlg_vec_tst is
end decoddisplay_vlg_vec_tst;
