library verilog;
use verilog.vl_types.all;
entity \trabalhofinalfinal__vlg_vec_tst\ is
end \trabalhofinalfinal__vlg_vec_tst\;
