library verilog;
use verilog.vl_types.all;
entity decoddisplay_vlg_check_tst is
    port(
        \OUT\           : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end decoddisplay_vlg_check_tst;
