library verilog;
use verilog.vl_types.all;
entity REG_2BYTES_vlg_vec_tst is
end REG_2BYTES_vlg_vec_tst;
